module Design_CHIP (
    I_clk, 
    I_rst, 
    O_done, 
    IO_F_IO_A, 
    O_F_CLE_A, 
    O_F_ALE_A, 
    O_F_REN_A, 
    O_F_WEN_A, 
    I_F_RB_A, 
    IO_F_IO_B, 
    O_F_CLE_B, 
    O_F_ALE_B, 
    O_F_REN_B, 
    O_F_WEN_B, 
    I_F_RB_B, 
    I_KEY
);
    
endmodule